module somador(
    input [31:0]a,
    output [31:0]b
);
assign b = a + 32'd4;


endmodule
