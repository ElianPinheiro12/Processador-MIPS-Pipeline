module somador(
    input [31:0]a,
    output [31:0]c
);
assign c = a + 32'd4;


endmodule